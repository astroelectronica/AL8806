.title KiCad schematic
.include "C:/AE/AL8806/_models/AL8806.spice.txt"
.include "C:/AE/AL8806/_models/C2012X7R2A104K125AE_p.mod"
.include "C:/AE/AL8806/_models/C3216C0G1H104K160AA_s.mod"
.include "C:/AE/AL8806/_models/DFLS230.spice.txt"
.include "C:/AE/AL8806/_models/PD_7345_744777115_15u.lib"
.include "C:/AE/AL8806/_models/XLamp-XBD-Spice.txt"
D4 /B2 /B3 XB-DGRN
D2 /A /B1 XB-DGRN
D3 /B1 /B2 XB-DGRN
XU4 /A /K C3216C0G1H104K160AA_s
D7 /B5 /K XB-DGRN
D5 /B3 /B4 XB-DGRN
D6 /B4 /B5 XB-DGRN
XU1 VCC 0 C2012X7R2A104K125AE_p
V1 /DIMM 0 PULSE(0 {VPUL} {DELAY} {TR} {TF} {DUTY} {CYCLE})
R1 /DIMM /CTRL {RCTRL}
D1 /SW VCC DI_DFLS230
XU2 /A 0 0 /CTRL /SW /SW 0 VCC AL8806
XU3 /SW /K PD_7345_744777115_15u
R2 VCC /A {RSET}
V2 VCC 0 {VSOURCE}
.end
